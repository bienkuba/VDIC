`timescale 1ns/1ps

package mult_pkg;
	`include "coverage.svh"
	`include "tpgen.svh"
	`include "scoreboard.svh"
	`include "testbench.svh"
endpackage : mult_pkg
	
	
	
	
	
	
